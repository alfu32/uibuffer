module tui_renderer
