module tui

pub fn test_color_create() {
}
