module tui
