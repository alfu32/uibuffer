module tui

////////////    Box Drawing[1]
////////////    Official Unicode Consortium code chart (PDF)
////////////            0	1	2	3	4	5	6	7	8	9	A	B	C	D	E	F
////////////    U+250x	─	━	│	┃	┄	┅	┆	┇	┈	┉	┊	┋	┌	┍	┎	┏
////////////    U+251x	┐	┑	┒	┓	└	┕	┖	┗	┘	┙	┚	┛	├	┝	┞	┟
////////////    U+252x	┠	┡	┢	┣	┤	┥	┦	┧	┨	┩	┪	┫	┬	┭	┮	┯
////////////    U+253x	┰	┱	┲	┳	┴	┵	┶	┷	┸	┹	┺	┻	┼	┽	┾	┿
////////////    U+254x	╀	╁	╂	╃	╄	╅	╆	╇	╈	╉	╊	╋	╌	╍	╎	╏
////////////    U+255x	═	║	╒	╓	╔	╕	╖	╗	╘	╙	╚	╛	╜	╝	╞	╟
////////////    U+256x	╠	╡	╢	╣	╤	╥	╦	╧	╨	╩	╪	╫	╬	╭	╮	╯
////////////    U+257x	╰	╱	╲	╳	╴	╵	╶	╷	╸	╹	╺	╻	╼	╽	╾	╿
////////////            0	1	2	3	4	5	6	7	8	9	A	B	C	D	E	F
////////////    U+258x	▀	▁	▂	▃	▄	▅	▆	▇	█	▉	▊	▋	▌	▍	▎	▏
////////////    U+259x	▐	░	▒	▓	▔	▕	▖	▗	▘	▙	▚	▛	▜	▝	▞	▟

////////////    ┌─────────┬─────────┐  ╔═════════╦═════════╗  ╓────────╥───────────╖  ╒══════════════════╤══════════════════════════╕
////////////    │         │         │  ║         ║         ║  ║        ║           ║  │                  │                          │
////////////    ├─────────┼─────────┤  ╠═════════╬═════════╣  ╟────────╫───────────╢  ╞══════════════════╪══════════════════════════╡
////////////    │         │         │  ║         ║         ║  ║        ║           ║  │                  │                          │
////////////    │         │         │  ║         ║         ║  ║        ║           ║  │                  │                          │
////////////    │         │         │  ║         ║         ║  ║        ║           ║  │                  │                          │
////////////    │         │         │  ║         ║         ║  ║        ║           ║  │                  │                          │
////////////    └─────────┴─────────┘  ╚═════════╩═════════╝  ╙────────╨───────────╜  ╘══════════════════╧══════════════════════════╛
////////////    ┌──────────────────────────────────────────────────────┐
////////////    │                   ╔═════════════╗ Some Text          │▒
////////////    │                   ║             ║                    │▒
////////////    │                   ║             ║                    │▒
////////////    │                   ╚═══════╦═════╝ in the box         │▒
////////////    │                           ║                          │▒
////////////    │                           ║                          │▒
////////////    ╞═════════╤═════════════════╩══════════════╤═══════════╡▒
////////////    │         │                                │           │▒
////////////    │         │                                │           │▒
////////////    │         │                                │           │▒
////////////    │         ├─────────────────┬──────────────┤           │▒
////////////    │         │                 │              │           │▒
////////////    │         │                 │              │           │▒
////////////    │         └─────────────────┴──────────────┘           │▒
////////////    │                                                      │▒
////////////    │                                                      │▒
////////////    └──────────────────────────────────────────────────────┘▒
////////////    ▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒▒

////////////        Code	Result	Description
////////////        U+2700	✀	Black safety scissors
////////////        U+2701	✁	Upper blade scissors
////////////        U+2702	✂	Black scissors
////////////        U+2703	✃	Lower blade scissors
////////////        U+2704	✄	White scissors
////////////        U+2705	✅	White heavy check mark
////////////        U+2706	✆	Telephone location sign
////////////        U+2707	✇	Tape drive
////////////        U+2708	✈	Airplane
////////////        U+2709	✉	Envelope
////////////        U+270A	✊	Raised fist
////////////        U+270B	✋	Raised hand
////////////        U+270C	✌	Victory hand
////////////        U+270D	✍	Writing hand
////////////        U+270E	✎	Lower right pencil
////////////        U+270F	✏	Pencil
////////////        U+2710	✐	Upper right pencil
////////////        U+2711	✑	White nib
////////////        U+2712	✒	Black nib
////////////        U+2713	✓	Check mark
////////////        U+2714	✔	Heavy check mark
////////////        U+2715	✕	Multiplication X
////////////        U+2716	✖	Heavy multiplication X
////////////        U+2717	✗	Ballot X
////////////        U+2718	✘	Heavy ballot X
////////////        U+2719	✙	Outlined Greek cross
////////////        U+271A	✚	Heavy Greek cross
////////////        U+271B	✛	Open center cross
////////////        U+271C	✜	Heavy open center cross
////////////        U+271D	✝	Latin cross
////////////        U+271E	✞	Shadowed white Latin cross
////////////        U+271F	✟	Outlined Latin cross
////////////        U+2720	✠	Maltese cross
////////////        U+2721	✡	Star of David
////////////        U+2722	✢	Four teardrop-spoked asterisk
////////////        U+2723	✣	Four balloon-spoked asterisk
////////////        U+2724	✤	Heavy four balloon-spoked asterisk
////////////        U+2725	✥	Four club-spoked asterisk
////////////        U+2726	✦	Black four-pointed star
////////////        U+2727	✧	White four-pointed star
////////////        U+2728	✨	Sparkles
////////////        U+2729	✩	Stress outlined white star
////////////        U+272A	✪	Circled white star
////////////        U+272B	✫	Open center black star
////////////        U+272C	✬	Black center white star
////////////        U+272D	✭	Outlined black star
////////////        U+272E	✮	Heavy outlined black star
////////////        U+272F	✯	Pinwheel star
////////////        U+2730	✰	Shadowed white star
////////////        U+2731	✱	Heavy asterisk
////////////        U+2732	✲	Open center asterisk
////////////        U+2733	✳	Eight spoked asterisk
////////////        U+2734	✴	Eight pointed black star
////////////        U+2735	✵	Eight pointed pinwheel star
////////////        U+2736	✶	Six pointed black star
////////////        U+2737	✷	Eight pointed rectilinear black star
////////////        U+2738	✸	Heavy eight pointed rectilinear black star
////////////        U+2739	✹	Twelve pointed black star
////////////        U+273A	✺	Sixteen pointed asterisk
////////////        U+273B	✻	Teardrop spoked asterisk
////////////        U+273C	✼	Open center teardrop spoked asterisk
////////////        U+273D	✽	Heavy teardrop spoked asterisk
////////////        U+273E	✾	Six petalled black and white florette
////////////        U+273F	✿	Black florette
////////////        U+2740	❀	White florette
////////////        U+2741	❁	Eight petalled outlined black florette
////////////        U+2742	❂	Circled open center eight pointed star
////////////        U+2743	❃	Heavy teardrop spoked pinwheel asterisk
////////////        U+2744	❄	Snowflake
////////////        U+2745	❅	Tight trifoliate snowflake
////////////        U+2746	❆	Heavy chevron snowflake
////////////        U+2747	❇	Sparkle
////////////        U+2748	❈	Heavy sparkle
////////////        U+2749	❉	Balloon spoked asterisk
////////////        U+274A	❊	Eight teardrop spoked propeller asterisk
////////////        U+274B	❋	Heavy eight teardrop spoked propeller asterisk
////////////        U+274C	❌	Cross mark
////////////        U+274D	❍	Shadowed white circle
////////////        U+274E	❎	Negative squared cross mark
////////////        U+274F	❏	Lower right drop-shadowed white square
////////////        U+2750	❐	Upper right drop-shadowed white square
////////////        U+2751	❑	Lower right shadowed white square
////////////        U+2752	❒	Upper right shadowed white square
////////////        U+2753	❓	Black question mark ornament
////////////        U+2754	❔	White question mark ornament
////////////        U+2755	❕	White exclamation mark ornament
////////////        U+2756	❖	Black diamond minus white X
////////////        U+2757	❗	Heavy exclamation mark symbol
////////////        U+2758	❘	Light vertical bar
////////////        U+2759	❙	Medium vertical bar
////////////        U+275A	❚	Heavy vertical bar
////////////        U+275B	❛	Heavy single turned comma quotation mark ornament
////////////        U+275C	❜	Heavy single comma quotation mark ornament
////////////        U+275D	❝	Heavy double turned comma quotation mark ornament
////////////        U+275E	❞	Heavy double comma quotation mark ornament
////////////        U+275F	❜	Heavy low single comma quotation mark ornament
////////////        U+2760	❞	Heavy low double comma quotation mark ornament
////////////        U+2761	❡	Curved stem paragraph sign ornament
////////////        U+2762	❢	Heavy exclamation mark ornament
////////////        U+2763	❣	Heavy heart exclamation mark ornament
////////////        U+2764	❤	Heavy black heart
////////////        U+2765	❥	Rotated heavy black heart bullet
////////////        U+2766	❦	Floral heart
////////////        U+2767	❧	Rotated floral heart bullet
////////////        U+2768	❨	Medium left parenthesis ornament
////////////        U+2769	❩	Medium right parenthesis ornament
////////////        U+276A	❪	Medium flattened left parenthesis ornament
////////////        U+276B	❫	Medium flattened right parenthesis ornament
////////////        U+276C	❬	Medium left-pointing angle bracket ornament
////////////        U+276D	❭	Medium right-pointing angle bracket ornament
////////////        U+276E	❮	Heavy left-pointing angle quotation mark ornament
////////////        U+276F	❯	Heavy right-pointing angle quotation mark ornament
////////////        U+2770	❰	Heavy left-pointing angle bracket ornament
////////////        U+2771	❱	Heavy right-pointing angle bracket ornament
////////////        U+2772	❲	Light left tortoise shell bracket ornament
////////////        U+2773	❳	Light right tortoise shell bracket ornament
////////////        U+2774	❴	Medium left curly bracket ornament
////////////        U+2775	❵	Medium left curly bracket ornament
////////////        U+2776	❶	Dingbat negative circled digit one
////////////        U+2777	❷	Dingbat negative circled digit two
////////////        U+2778	❸	Dingbat negative circled digit three
////////////        U+2779	❹	Dingbat negative circled digit four
////////////        U+277A	❺	Dingbat negative circled digit five
////////////        U+277B	❻	Dingbat negative circled digit six
////////////        U+277C	❼	Dingbat negative circled digit seven
////////////        U+277D	❽	Dingbat negative circled digit eight
////////////        U+277E	❾	Dingbat negative circled digit nine
////////////        U+277F	❿	Dingbat negative circled digit ten
////////////        U+2780	➀	Dingbat circled sans-serif digit one
////////////        U+2781	➁	Dingbat circled sans-serif digit two
////////////        U+2782	➂	Dingbat circled sans-serif digit three
////////////        U+2783	➃	Dingbat circled sans-serif digit four
////////////        U+2784	➄	Dingbat circled sans-serif digit five
////////////        U+2785	➅	Dingbat circled sans-serif digit six
////////////        U+2786	➆	Dingbat circled sans-serif digit seven
////////////        U+2787	➇	Dingbat circled sans-serif digit eight
////////////        U+2788	➈	Dingbat circled sans-serif digit nine
////////////        U+2789	➉	Dingbat circled sans-serif digit ten
////////////        U+278A	➊	Dingbat negative circled sans-serif digit one
////////////        U+278B	➋	Dingbat negative circled sans-serif digit two
////////////        U+278C	➌	Dingbat negative circled sans-serif digit three
////////////        U+278D	➍	Dingbat negative circled sans-serif digit four
////////////        U+278E	➎	Dingbat negative circled sans-serif digit five
////////////        U+278F	➏	Dingbat negative circled sans-serif digit six
////////////        U+2790	➐	Dingbat negative circled sans-serif digit seven
////////////        U+2791	➑	Dingbat negative circled sans-serif digit eight
////////////        U+2792	➒	Dingbat negative circled sans-serif digit nine
////////////        U+2793	➓	Dingbat negative circled sans-serif digit ten
////////////        U+2794	➔	Heavy wide-headed rightward arrow
////////////        U+2795	➕	Heavy plus sign
////////////        U+2796	➖	Heavy minus sign
////////////        U+2797	➗	Heavy division sign
////////////        U+2798	➘	Heavy south east arrow
////////////        U+2799	➙	Heavy rightward arrow
////////////        U+279A	➚	Heavy north east arrow
////////////        U+279B	➛	Drafting point rightward arrow
////////////        U+279C	➜	Heavy round-tipped rightward arrow
////////////        U+279D	➝	Triangle-headed rightward arrow
////////////        U+279E	➞	Heavy triangle-headed rightward arrow
////////////        U+279F	➟	Dashed triangle-headed rightward arrow
////////////        U+27A0	➠	Heavy dashed triangle-headed rightward arrow
////////////        U+27A1	➡	Black rightward arrow
////////////        U+27A2	➢	Three-D top-lighted rightward arrowhead
////////////        U+27A3	➣	Three-D bottom-lighted rightward arrowhead
////////////        U+27A4	➤	Black rightward arrowhead
////////////        U+27A5	➥	Heavy black curved downward and rightward arrow
////////////        U+27A6	➦	Heavy black curved upward and rightward arrow
////////////        U+27A7	➧	Squat black rightward arrow
////////////        U+27A8	➨	Heavy concave-pointed black rightward arrow
////////////        U+27A9	➩	Right-shaded white rightward arrow
////////////        U+27AA	➪	Left-shaded white rightward arrow
////////////        U+27AB	➫	Back-tilted shadowed white rightward arrow
////////////        U+27AC	➬	Front-tilted shadowed white rightward arrow
////////////        U+27AD	➭	Heavy lower right-shadowed white rightward arrow
////////////        U+27AE	➮	Heavy upper right-shadowed white rightward arrow
////////////        U+27AF	➯	Notched lower right-shadowed white rightward arrow
////////////        U+27B0	➰	Curly loop
////////////        U+27B1	➱	Notched upper right-shadowed white rightward arrow
////////////        U+27B2	➲	Circled heavy white rightward arrow
////////////        U+27B3	➳	White-feathered rightward arrow
////////////        U+27B4	➴	Black-feathered south east arrow
////////////        U+27B5	➵	Black-feathered rightward arrow
////////////        U+27B6	➶	Black-feathered north east arrow
////////////        U+27B7	➷	Heavy black-feathered south east arrow
////////////        U+27B8	➸	Heavy black-feathered rightward arrow
////////////        U+27B9	➹	Heavy black-feathered north east arrow
////////////        U+27BA	➺	Teardrop-barbed rightward arrow
////////////        U+27BB	➻	Heavy teardrop-shanked rightward arrow
////////////        U+27BC	➼	Wedge-tailed rightward arrow
////////////        U+27BD	➽	Heavy wedge-tailed rightward arrow
////////////        U+27BE	➾	Open-outlined rightward arrow
////////////        U+27BF	➿	Double curly loop
