module tui_renderer

pub fn test_color_create() {
}
